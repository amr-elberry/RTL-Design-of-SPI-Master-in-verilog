/****************************************time scale*************************************/
`timescale 1ns/1ps
/***************************************************************************************/


/***********************************declara tb signal***********************************/
module clk_div_tb (
	input reg clk_tb,rst_tb,valid_tb,
	output wire leading_edge_tb,trailing_edge_tb,clk_div_tb
	);
/***************************************************************************************/


/****************************DUT instantiation******************************************/
DUT clk_div_tb(
.clk(clk_tb),
.clk_div(clk_div_tb),
.rst(rst_tb).
.valid(valid_tb)
.leading_edge(leading_edge_tb),
.trailing_edge(trailing_edge_tb));


/***************************************************************************************/

/*****************************tasks****************************************************/



/**************************************************************************************/

/********************************** intial block **************************************/
initial
begin
	$dumpvars
	$dumpfile(clk_TB.vcd)
	
end

/**************************************************************************************/